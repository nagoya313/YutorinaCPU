`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

`include "bus.h"

module bus(input wire clock, input wire reset,
           output wire [`YutorinaWordDataBus] master_read_data,
           output wire master_ready_,
           input wire master0_request_, 
           input wire [`YutorinaWordAddressBus] master0_address,
           input wire master0_address_strobe_,
           input wire master0_read_write,
           input wire [`YutorinaWordDataBus] master0_write_data,
           output wire master0_grant_,
           input wire master1_request_, 
           input wire [`YutorinaWordAddressBus] master1_address,
           input wire master1_address_strobe_,
           input wire master1_read_write,
           input wire [`YutorinaWordDataBus] master1_write_data,
           output wire master1_grant_,
           input wire master2_request_, 
           input wire [`YutorinaWordAddressBus] master2_address,
           input wire master2_address_strobe_,
           input wire master2_read_write,
           input wire [`YutorinaWordDataBus] master2_write_data,
           output wire master2_grant_,
           input wire master3_request_, 
           input wire [`YutorinaWordAddressBus] master3_address,
           input wire master3_address_strobe_,
           input wire master3_read_write,
           input wire [`YutorinaWordDataBus] master3_write_data,
           output wire master3_grant_,
           output wire [`YutorinaWordAddressBus] slave_address,
           output wire slave_address_strobe_,
           output wire slave_read_write,
           output wire [`YutorinaWordDataBus] slave_write_data,
           input wire [`YutorinaWordDataBus] slave0_read_data,
           input wire slave0_ready_, output wire slave0_chip_select_,
           input wire [`YutorinaWordDataBus] slave1_read_data,
           input wire slave1_ready_, output wire slave1_chip_select_,
           input wire [`YutorinaWordDataBus] slave2_read_data,
           input wire slave2_ready_, output wire slave2_chip_select_,
           input wire [`YutorinaWordDataBus] slave3_read_data,
           input wire slave3_ready_, output wire slave3_chip_select_,
           input wire [`YutorinaWordDataBus] slave4_read_data,
           input wire slave4_ready_, output wire slave4_chip_select_,
           input wire [`YutorinaWordDataBus] slave5_read_data,
           input wire slave5_ready_, output wire slave5_chip_select_,
           input wire [`YutorinaWordDataBus] slave6_read_data,
           input wire slave6_ready_, output wire slave6_chip_select_,
           input wire [`YutorinaWordDataBus] slave7_read_data,
           input wire slave7_ready_, output wire slave7_chip_select_);
  bus_arbiter bus_arbiter(.clock (clock), .reset (reset),
                          .master0_request_ (master0_request_),
                          .master0_grant_ (master0_grant_),
                          .master1_request_ (master1_request_),
                          .master1_grant_ (master1_grant_),
                          .master2_request_ (master2_request_),
                          .master2_grant_ (master2_grant_),
                          .master3_request_ (master3_request_),
                          .master3_grant_ (master3_grant_));
  bus_master_multiplexer bus_master_multiplexer(
    .master0_address (master0_address), 
    .master0_address_strobe_ (master0_address_strobe_),
    .master0_read_write (master0_read_write),
    .master0_write_data (master0_write_data),
    .master0_grant_ (master0_grant_),
    .master1_address (master1_address), 
    .master1_address_strobe_ (master1_address_strobe_),
    .master1_read_write (master1_read_write),
    .master1_write_data (master1_write_data),
    .master1_grant_ (master1_grant_),
    .master2_address (master1_address), 
    .master2_address_strobe_ (master2_address_strobe_),
    .master2_read_write (master2_read_write),
    .master2_write_data (master2_write_data),
    .master2_grant_ (master2_grant_),
    .master3_address (master3_address), 
    .master3_address_strobe_ (master3_address_strobe_),
    .master3_read_write (master3_read_write),
    .master3_write_data (master3_write_data),
    .master3_grant_ (master3_grant_),
    .slave_address (slave_address),
    .slave_address_strobe_ (slave_address_strobe_),
    .slave_read_write (slave_read_write),
    .slave_write_data (slave_write_data));
  bus_address_decoder bus_address_decoder(
    .slave_address (slave_address),
    .slave0_chip_select_ (slave0_chip_select_),
    .slave1_chip_select_ (slave1_chip_select_),
    .slave2_chip_select_ (slave2_chip_select_),
    .slave3_chip_select_ (slave3_chip_select_),
    .slave4_chip_select_ (slave4_chip_select_),
    .slave5_chip_select_ (slave5_chip_select_),
    .slave6_chip_select_ (slave6_chip_select_),
    .slave7_chip_select_ (slave7_chip_select_));
  bus_slave_multiplexer bus_slave_multiplexer(
    .slave0_chip_select_ (slave0_chip_select_), 
    .slave1_chip_select_ (slave1_chip_select_),
    .slave2_chip_select_ (slave2_chip_select_),
    .slave3_chip_select_ (slave3_chip_select_),
    .slave4_chip_select_ (slave4_chip_select_),
    .slave5_chip_select_ (slave5_chip_select_),
    .slave6_chip_select_ (slave6_chip_select_),
    .slave7_chip_select_ (slave7_chip_select_),
    .slave0_read_data (slave0_read_data), .slave0_ready_ (slave0_ready_),
    .slave1_read_data (slave1_read_data), .slave1_ready_ (slave1_ready_),
    .slave2_read_data (slave2_read_data), .slave2_ready_ (slave2_ready_),
    .slave3_read_data (slave3_read_data), .slave3_ready_ (slave3_ready_),
    .slave4_read_data (slave4_read_data), .slave4_ready_ (slave4_ready_),
    .slave5_read_data (slave5_read_data), .slave5_ready_ (slave5_ready_),
    .slave6_read_data (slave6_read_data), .slave6_ready_ (slave6_ready_),
    .slave7_read_data (slave7_read_data), .slave7_ready_ (slave7_ready_),
    .master_read_data (master_read_data), .master_ready_(master_ready_));
endmodule
