`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

`timescale 1ns/1ps

module yutorina_clk_gen(
  input wire clk_ref, input wire rst_sw,
  output wire clk, output wire clk_, output wire chip_rst);
  wire locked;
  wire dcm_rst;
  assign dcm_rst = (rst_sw == `RESET_ENABLE) ? `ENABLE : `DISABLE;
  assign chip_rst = (rst_sw == `RESET_ENABLE) || (locked == `DISABLE) ?
                     `ENABLE : `DISABLE;
  // ざいりんくすの何か
  x_s3e_dcm x_s3e_dcm(.CLKIN_IN (clk_ref), .RST_IN (dcm_rst),
                      .CLK0_OUT (clk), .CLK180_OUT (clk_),
                      .LOCKED_OUT (locked));
endmodule
